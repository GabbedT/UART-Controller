import UART_pkg::*;

module interrupt_arbiter (
  input  logic       clk_i,
  input  logic       rst_n_i,
  input  logic       rx_dsm_i,

  /* Interrupt cause */
  input  logic       rx_rdy_i,
  input  logic       tx_done_i,
  input  logic       cfg_error_i,
  input  logic       parity_error_i,
  input  logic       frame_error_i,
  input  logic       overrun_error_i,
  input  logic       rx_fifo_full_i,
  input  logic       config_req_slv_i,

  /* Enable interrupt */
  input  logic       overrun_error_en_i,
  input  logic       frame_error_en_i,
  input  logic       parity_error_en_i,
  input  logic       rx_rdy_en_i,

  /* Interrupt clear */
  input  logic       int_ackn_i,
  input  logic       config_ackn_i,
  input  logic       read_rx_data_i,
  input  logic       rx_fifo_empty_i,

  output logic [2:0] interrupt_vector_o,
  output logic       irq_n_o
);

  /* Next and current state */
  localparam NXT = 1;
  localparam CRT = 0;

  typedef struct packed {
    /* Valid when = 0 */
    logic       valid_n;
    logic [2:0] vector;
  } interrupt_t;


//--------------------//
//  ENABLE INTERRUPT  //
//--------------------//

  logic overrun_error, parity_error, frame_error, rx_rdy;

  assign overrun_error = overrun_error_i & overrun_error_en_i;
  assign parity_error = parity_error_i & parity_error_en_i;
  assign frame_error = frame_error_i & frame_error_en_i;
  assign rx_rdy = rx_rdy_i & rx_rdy_en_i;


//-------------------//
//  PRIORITY 1 FIFO  //
//-------------------//

  logic prio1_fifo_write;

  assign prio1_fifo_write = cfg_error_i | parity_error | frame_error | overrun_error;

  /* FIFO interface assignment */
  sync_fifo_interface #(4) fifo_prio1_if(clk_i);

  assign fifo_prio1_if.write_i = prio1_fifo_write;
  assign fifo_prio1_if.rst_n_i = rst_n_i;
  assign fifo_prio1_if.wr_data_i = {cfg_error_i, overrun_error, frame_error, parity_error};


  /* FIFO buffer instantiation in FWFT mode */
  sync_FIFO_buffer #(4, 1) priority1_fifo (fifo_prio1_if);

  logic [3:0] prio1_data_read[NXT:CRT];

      always_ff @(posedge clk_i) begin 
        if (!rst_n_i) begin 
          prio1_data_read[CRT] <= 2'b0;
        end else begin 
          prio1_data_read[CRT] <= prio1_data_read[NXT];
        end
      end

  /* Vector generated by first priority interrupt */
  logic [2:0] prio1_int_vector;

      always_comb begin : prio1_vector_gen
        /* Internal priority:
         * -------------------------------------------------------
         *    - CONFIGURATION ERROR
         *    - OVERRUN ERROR
         *    - FRAME ERROR 
         *    - PARITY ERROR
         */
        casez (prio1_data_read[CRT])
          4'b1???: prio1_int_vector = {1'b0, INT_CONFIG_FAIL};
          4'b01??: prio1_int_vector = {1'b0, INT_OVERRUN};
          4'b001?: prio1_int_vector = {1'b0, INT_FRAME};
          4'b0001: prio1_int_vector = {1'b0, INT_PARITY};
          default: prio1_int_vector = {1'b1, 3'b000};
        endcase
      end : prio1_vector_gen


//-------------------//
//  PRIORITY 2 FIFO  //
//-------------------//

  logic prio2_fifo_write;

  assign prio2_fifo_write = rx_fifo_full_i | config_req_slv_i;

  /* FIFO interface assignment */
  sync_fifo_interface #(2) fifo_prio2_if(clk_i);

  assign fifo_prio2_if.write_i = prio2_fifo_write;
  assign fifo_prio2_if.rst_n_i = rst_n_i;
  assign fifo_prio2_if.wr_data_i = {rx_fifo_full_i, config_req_slv_i};

  /* FIFO buffer instantiation in FWFT mode */
  sync_FIFO_buffer #(4, 1) priority2_fifo (fifo_prio2_if);

  logic [1:0] prio2_data_read[NXT:CRT];

      always_ff @(posedge clk_i) begin 
        if (!rst_n_i) begin 
          prio2_data_read[CRT] <= 2'b0;
        end else begin 
          prio2_data_read[CRT] <= prio2_data_read[NXT];
        end
      end

  /* Vector generated by second priority interrupt */
  interrupt_t prio2_int_vector;

      always_comb begin : prio2_vector_gen
        /* Internal priority:
         * -------------------------------------------------------
         *    - RECEIVER FIFO FULL
         *    - REQUESTED CONFIGURATION
         */
        casez (prio2_data_read[CRT])
          2'b1?:   prio2_int_vector = {1'b0, INT_RX_FULL};
          2'b01:   prio2_int_vector = {1'b0, INT_CONFIG_REQ};
          default: prio2_int_vector = {1'b1, 3'b000};
        endcase
      end : prio2_vector_gen


//-------------------//
//  PRIORITY 3 FIFO  //
//-------------------//

  logic prio3_fifo_write;

  assign prio3_fifo_write = tx_done_i | rx_rdy;

  sync_fifo_interface #(2) fifo_prio3_if(clk_i);

  assign fifo_prio3_if.write_i = prio3_fifo_write;   
  assign fifo_prio3_if.rst_n_i = rst_n_i;         
  assign fifo_prio3_if.wr_data_i = {rx_rdy, tx_done_i};

  /* FIFO buffer instantiation in FWFT mode */
  sync_FIFO_buffer #(4, 1) priority3_fifo (fifo_prio3_if);

  logic [1:0] prio3_data_read[NXT:CRT];

      always_ff @(posedge clk_i) begin 
        if (!rst_n_i) begin 
          prio3_data_read[CRT] <= 2'b0;
        end else begin 
          prio3_data_read[CRT] <= prio3_data_read[NXT];
        end
      end

  /* Vector generated by third priority interrupt */
  interrupt_t prio3_int_vector;

      always_comb begin : prio3_vector_gen
        /* Internal priority:
         * -------------------------------------------------------
         *    - DATA RECEIVED READY
         *    - TRANSMISSION DONE
         */        
        casez (prio3_data_read[CRT])
          2'b1?:   prio3_int_vector = {1'b0, INT_RXD_RDY};
          2'b01:   prio3_int_vector = {1'b0, INT_TX_DONE};
          default: prio3_int_vector = {1'b1, 3'b000};
        endcase
      end : prio3_vector_gen


//---------------------//
//  PRIORITY SELECTOR  // 
//---------------------//

  logic PRIORITY_1 = 3'b??1;
  logic PRIORITY_2 = 3'b?10;
  logic PRIORITY_3 = 3'b100;

  /* One hot selector */
  logic [2:0] priority_select;

  assign priority_select[0] = !fifo_prio1_if.empty_o;
  assign priority_select[1] = !fifo_prio2_if.empty_o;
  assign priority_select[2] = !fifo_prio3_if.empty_o;

  interrupt_t interrupt; 

      /* Select the interrupt with highest priority */
      always_comb begin 
        casez (priority_select)
          PRIORITY_1: interrupt = prio1_int_vector;
          PRIORITY_2: interrupt = prio2_int_vector;
          PRIORITY_3: interrupt = prio3_int_vector;
          default:    interrupt = {1'b1, 3'b000};
        endcase
      end

  assign interrupt_vector_o = interrupt.vector;

  logic irq_n;

      always_ff @(posedge clk_i) begin 
        if (!rst_n_i) begin 
          irq_n_o <= 1'b1;
        end else begin 
          irq_n_o <= irq_n;
        end
      end

  typedef enum logic [1:0] {
    IDLE,
    /* Retrieve interrupt vector */
    READ_VECTOR,
    /* Wait interrupt to be cleared */
    WAIT_ACKN,
    /* IRQ should stay low for at least 1 clock cycle */
    CLEAR,
  } arbiter_fsm_e;


      always_comb begin : acknowledge_logic
        /* Default values */
        fifo_prio1_if.read_i = priority_select[0];
        fifo_prio2_if.read_i = priority_select[1];
        fifo_prio3_if.read_i = priority_select[2];
        prio1_data_read[NXT] = fifo_prio1_if.rd_data_o;
        prio2_data_read[NXT] = fifo_prio2_if.rd_data_o;
        prio3_data_read[NXT] = fifo_prio3_if.rd_data_o;
        irq_n = interrupt.valid_n;

        /* If the interrupt get acknowlege, before getting the new
         * interrupt bundle (reading the fifo to get the next 
         * interrupt) check if in the same bundle there's another
         * interrupt to acknowledge. If there's one, clear the 
         * preceeding one and process the next one. */
        if (!interrupt.valid_n) begin
          case (interrupt.vector)
            INT_TX_DONE: begin 
              fifo_prio3_if.read_i = int_ackn_i & (!prio3_data_read[CRT][1]);
              irq_n = fifo_prio3_if.read_i;

              if (!prio3_data_read[CRT][1]) begin
                prio3_data_read[NXT] = fifo_prio3_if.rd_data_o;
              end else begin 
                prio3_data_read[NXT] = {prio3_data_read[CRT][1], 1'b0};
              end
            end   

            INT_CONFIG_FAIL: begin  
              fifo_prio1_if.read_i = int_ackn_i & (prio1_data_read[CRT][2:0] == 3'b0);
              irq_n = !fifo_prio1_if.read_i;

              if (prio1_data_read[CRT][2:0] == 3'b0) begin 
                prio1_data_read[NXT] = fifo_prio1_if.rd_data_o;
              end else begin 
                prio1_data_read[NXT] = {1'b0, prio1_data_read[CRT][2:0]};
              end
            end 

            /* Those 3 interrupt require a data read, that will clear 
            * the other ones too if there are multiple interrupt in
            * a transaction. */
            INT_OVERRUN: begin 
              fifo_prio1_if.read_i = read_rx_data_i;
              irq_n = !fifo_prio1_if.read_i;
            end

            INT_FRAME: begin 
              fifo_prio1_if.read_i = read_rx_data_i;
              irq_n = !fifo_prio1_if.read_i;
            end

            INT_PARITY: begin 
              fifo_prio1_if.read_i = read_rx_data_i;
              irq_n = !fifo_prio1_if.read_i;
            end

            INT_RXD_RDY: begin  
              fifo_prio3_if.read_i = ((rx_dsm_i) ? rx_fifo_empty_i : read_rx_data_i) & (!prio3_data_read[CRT][0]);
              irq_n = !fifo_prio3_if.read_i;

              if (!prio3_data_read[CRT][0]) begin
                prio3_data_read[NXT] = fifo_prio3_if.rd_data_o;
              end else begin 
                prio3_data_read[NXT] = {1'b0, prio3_data_read[CRT][0]};
              end
            end

            INT_RX_FULL: begin 
              fifo_prio2_if.read_i = ((rx_dsm_i) ? rx_fifo_empty_i : read_rx_data_i) & (!prio2_data_read[CRT][0]);
              irq_n = !fifo_prio2_if.read_i;

              if (!prio2_data_read[CRT][0]) begin
                prio2_data_read[NXT] = fifo_prio2_if.rd_data_o;
              end else begin 
                prio2_data_read[NXT] = {1'b0, prio2_data_read[CRT][0]};
              end            
            end

            INT_CONFIG_REQ: begin 
              fifo_prio2_if.read_i = config_ackn_i & (!prio2_data_read[CRT][1]);
              irq_n = !fifo_prio2_if.read_i;

              if (!prio2_data_read[CRT][1]) begin
                prio2_data_read[NXT] = fifo_prio2_if.rd_data_o;
              end else begin 
                prio2_data_read[NXT] = {prio2_data_read[CRT][1], 1'b0};
              end  
            end
          endcase
        end
      end : acknowledge_logic

endmodule